.SUBCKT  L_744834101_1m  1  2  3  4 PARAMS:
+  L1=200.14u
+  L2=200.53u
+  L3=254.10u
+  L4=250.1u
+  L5=10n
+  C1=18000.06f
+  C2=540.02f
+  Rs1=1856.63
+  Rs2=1278.77
+  Rs3=1496.33
+  Rs4=18000
+  Rs5=1636.33
+  R2=7
+  dL3=380e-009
+  dC3=6.5e-012
+  dL4=13.51e-009
+  dC4=7.63e-012
+  dR3=0.48
+  dR4=3550
+  dR5=0.78
+  dR6=466
+  Rdc=8m
+  ck=2pF
R_R9  N12325  3  {R2}
R_R8  N13265  N13287  {Rs4} 
Kn_K6 L_L11 L_L12 0.9999
Kn_K7 L_L11 L_L13 0.9999
Kn_K8 L_L11 L_L14 0.9999
Kn_K9 L_L12 L_L13 0.9999
Kn_K10 L_L12 L_L14 0.9999
Kn_K11 L_L13 L_L14 0.9999
R_R3  N12571  N12583  {Rs3}
R_R10  N13777  4  {R2}
C_C10  N13029  N12821  {ck}
R_R20  N13215  N13229  {dR4}
L_L11  N12821  N12295  {dL4}
R_R17  N12267  N12273  {dR3}
L_L8  N13265  N13287  {L4}
R_R7  N13287  N13305  {Rs3}
L_L9  N12295  N12307  {L5}
Kn_K4  L_L7  L_L8  1
R_R2  N12583  N12599  {Rs2}
Kn_K5  L_L9  L_L10  1
R_R16  N13229  N13249  {dR6}
Kn_K12 L_L15 L_L16 0.9999
Kn_K13 L_L15 L_L17 0.9999
Kn_K14 L_L15 L_L18 0.9999
Kn_K15 L_L16 L_L17 0.9999
Kn_K16 L_L16 L_L18 0.9999
Kn_K17 L_L17 L_L18 0.9999
C_C5  N12273  N12289  {dC4}
L_L6  N13287  N13305  {L3}
L_L7  N12307  N12571  {L4}
R_R6  N13305  N13319  {Rs2}
R_R21  1  N12257  {Rdc}
Kn_K3  L_L5  L_L6  1
L_L16  N12257  N12799  {dL3}
C_C8  N13215  N13741  {dC3}
L_L18  N13023  N13215  {dL3}
R_R1  N12599  3  {Rs1}
R_R13  N12289  N12295  {dR5}
L_L4  N13305  N13319  {L2}
L_L5  N12571  N12583  {L3}
R_R15  N13755  N13249  {dR5}
R_R5  N13319  4  {Rs1}
R_R18  N12257  N12273  {dR4}
Kn_K2  L_L3  L_L4  1
R_R19  N13741  N13229  {dR3}
L_L15  N12799  N12273  {dL3}
L_L17  N13229  N13023  {dL3}
L_L3  N12583  N12599  {L2}
R_R11  N12295  N12307  {Rs5}
L_L2  N13319  4  {L1}
C_C4  N13249  N13265  {C2}
L_L10  N13249  N13265  {L5}
Kn_K1  L_L1  L_L2  1
R_R14  N12273  N12295  {dR6}
C_C6  N13229  N13755  {dC4}
L_L12  N12273  N12821  {dL4}
L_L14  N13029  N13229  {dL4}
L_L1  N12599  3  {L1}
C_C1  N12307  N12325  {C1}
R_R12  N13249  N13265  {Rs5}
C_C2  N13265  N13777  {C1}
R_R22  2  N13215  {Rdc}
C_C9  N13023  N12799  {ck}
R_R4  N12307  N12571  {Rs4}
C_C3  N12295  N12307  {C2}
L_L13  N13249  N13029  {dL4}
C_C7  N12257  N12267  {dC3}
.ends  L_744834101_1m
******